module ControlUnit(opcode, ALU, REG, immediate, memWrite, memOut, );
  
