module InstMem(address, clk, out);
  input[15:0] address;
  input clk;
  output reg[31:0] out;
  integer firstclock = 0;

  reg[31:0] mem[16:0];
  
  always@(posedge clk)
  begin
	if(firstclock == 0)
	begin
		// instruções
		
		mem[0] = 32'b01011000000000010000000000000000;
		mem[1] = 32'b01011100000000010000000000000000;
		mem[2] = 32'b00000100001000000001000000000000;
		mem[3] = 32'b01000000001000100001100000000000;
		mem[4] = 32'b01011100000000110000000000000000;
		mem[5] = 32'b01001000000000110000000000000001;
		mem[6] = 32'b01100100000001000000000000000011;
		mem[7] = 32'b01100100000001000000000000000100;
		mem[8] = 32'b01110100000001000000000000000000;
		mem[9] = 32'b01100000000001010000000000000000;
		mem[10] = 32'b01011100000001010000000000000000;
		mem[11] = 32'b00110000101000000010100001000000;
		mem[12] = 32'b01011100000001010000000000000000;
		mem[13] = 32'b00000000000000000000000000000000;
		mem[14] = 32'b01001100000000000000000000000000;

 		
		firstclock <= 1;
	end
  end

  

  always@(address)
  begin
    out = mem[address];
  end

endmodule
